
module execute(
  input clk,
  input reset,

  // from decode to execute
  input         decode_valid, 
  output        decode_retry, 
  input  [31:0] decode_insn, 
  input  [63:0] decode_pc,
  input  [63:0] decode_sign_ext, 
  input  [63:0] decode_src1, 
  input  [63:0] decode_src2,

  // from execute to fetch
  output           execute_valid,
  input            execute_retry, // ALWAYS FALSE from fetch
  output  [63-1:0] execute_pc,

  // from execute to decode
  output        dest_valid,
  input         dest_retry, // ALWAYS FALSE from decode
  output [4:0]  dest_rd,
  output        dest_long,
  output [63:0] dest_data,
  output        dest_clear, // Just clear dependence, do not write to register

  // dcache interface (from execute to testbench)
  output [63:0] dcache_req_addr,  // load or store address computed at execute
  output [63:0] dcache_req_data, // data just for the store going to from exe to testbench
  output [3:0]  dcache_req_op,  // RVMOP_*
  output [4:0]  dcache_req_rd,  // destination register for the load
  output        dcache_req_valid,
  input         dcache_req_retry
);


  localparam  LOAD      = 7'b0000011;
  localparam  OP_IMM    = 7'b0010011;
  localparam  OP_IMM_32 = 7'b0011011;
  localparam  STORE     = 7'b0100011;
  localparam  OP        = 7'b0110011;
  localparam  OP_32     = 7'b0111011;
  localparam  BRANCH    = 7'b1100011;
  localparam  JALR      = 7'b1100111;


// LAB4 Main new thing:
//
// -Handle back to back instruction (dependences) (last_dest and last_reg...)
//
// -Compute LD/ST operations and send to testbench
//
// -PC+4 is generated by fetch, but checked here
//
// -Discard instructions that got incorrectly fetched. Discard instructions until the fix PC
// gets to execute.
//
// -When discarding instructions, some instructions can be stalled at decode
// due to wait for a load. Clear pending from execute to decode (no retry
// allowed). Set the dest_clear and ingore the dest_data when a load that
// needs to be flushed reaches execute


//flop_r #(.Reset_Value(1)) f_valid ( .d(decode_valid), .q(execute_valid),.*);
//assign decode_retry = 1'b0;
//flop f_retry ( .d(execute_retry), .q(decode_retry), .*);
wire [6:0] operation;
assign operation = decode_insn[6:0];


wire [63:0] pc;

//flop #(.Bits(64)) delay_pc ( .d(decode_pc), .q(pc), .*);
//flop_er #(.Bits(64),.Reset_Value(64'b0)) f_pc ( .d(decode_pc+4), .q(pc), .we(decode_valid), .*);

wire [4:0] rs1;
wire [4:0] rs2;
assign rs2 = decode_insn[24:20];
assign rs1 = decode_insn[19:15];

//remember last 2 rd
assign current_rd = dest_rd; 
wire [4:0] current_rd;
wire [4:0] last_rd;
wire [4:0] twolast_rd;
wire [4:0] threelast_rd;

wire last_valid;
wire twolast_valid;
wire threelast_valid;

//remember last 2 rd_data
assign current_data = dest_data;
wire [63:0] current_data;
wire [63:0] last_data;
wire [63:0] twolast_data;
wire [63:0] threelast_data;

fflop #(.Size(64+5)) rd_mem1 ( 
  .din({current_rd, current_data}), 
  .dinValid(dest_valid),
  .dinRetry(),
  
  .q({last_rd, last_data}),
  .qValid(last_valid),
  .qRetry(dcache_req_retry), 
  .*);
fflop #(.Size(64+5)) rd_mem2 ( 
  .din({last_rd, last_data}),  
  .dinValid(last_valid),
  .dinRetry(),

  .q({twolast_rd,twolast_data}),
  .qValid(twolast_valid),
  .qRetry(dcache_req_retry), 
 
  .*);
fflop #(.Size(64+5)) rd_mem3 ( 
  .din({twolast_rd, twolast_data}),  
  .dinValid(twolast_valid),
  .dinRetry(),

  .q({threelast_rd, threelast_data}), 
  .qValid(threelast_valid),
  .qRetry(dcache_req_retry), 
 
  .*);
/*
fflop #(.Size(64)) data_mem1 ( 
  .din(current_data),  
  .dinValid(dest_valid),
  .dinRetry(),

  .q(last_data), 
  .qValid(last_valid),
  .qRetry(dcache_req_retry), 
 
  .*);
fflop #(.Size(64)) data_mem2 ( 
  .din(last_data),  
  .dinValid(last_valid),
  .dinRetry(),

  .q(twolast_data), 
  .qValid(twolast_valid),
  .qRetry(dcache_req_retry), 
 
  .*);
fflop #(.Size(64)) data_mem3 ( 
  .din(twolast_data),  
  .dinValid(twolast_valid),
  .dinRetry(),

  .q(threelast_data), 
  .qValid(threelast_valid),
  .qRetry(dcache_req_retry), 
 
  .*);
*/
/*
reg [4:0] current_rd;
reg [4:0] last_rd;
reg [4:0] twolast_rd;
reg [4:0] threelast_rd;

reg [63:0] current_data;
reg [63:0] last_data;
reg [63:0] twolast_data;
reg [63:0] threelast_data;
always @(*) begin
  if(dest_valid) begin
    current_rd = dest_rd;
    current_data = dest_data;
  end
end
*/

reg [63:0]  rs1_data;
reg [63:0]  rs2_data;

always @ (*) begin
  if(operation == OP ||operation == OP_IMM ||operation == OP_IMM_32 ||operation == OP_32 ||operation == BRANCH ||operation == JALR ||operation == LOAD ||operation == STORE) begin
    if(rs1 == current_rd && dest_valid) begin
      rs1_data = current_data;
    end else if(rs1 == last_rd && last_valid) begin
      rs1_data = last_data;
    end else if(rs1 == twolast_rd && twolast_valid) begin
      rs1_data = twolast_data;
    end else if(rs1 == threelast_rd && threelast_valid) begin
      rs1_data = threelast_data;
    end else begin 
      $display("1NONE");
      rs1_data = decode_src1;
    end
  end
  if(operation == OP || operation == OP_32 || operation == BRANCH || operation == STORE) begin
    if(rs2 == current_rd &&dest_valid) begin
      rs2_data = current_data;
    end else if(rs2 == last_rd && last_valid) begin
      rs2_data = last_data;
    end else if(rs2 == twolast_rd && twolast_valid) begin
      rs2_data = twolast_data;
    end else if(rs2 == threelast_rd && threelast_valid) begin
      rs2_data = threelast_data;
    end else begin
      $display("2NONE");
      rs2_data = decode_src2;
    end
  end 

 // $display("reg = %d, CURRENT_RD = %d", current_rd,current_data);
 // $display("reg = %d, LAST_RD = %d", last_rd,last_data);
 // $display("reg = %d, TWOLAST_RD = %d", twolast_rd,twolast_data);
 // $display("reg = %d, THREELAST_RD = %d", threelast_rd,threelast_data);
 // $display("%d USED1 = %d, %d USED2 = %d", rs1, rs1_data, rs2, rs2_data);
end

// instantiate ALU here
alu a (
  .clk(clk),
  .reset(reset),

  // All the inputs come from decode stage
  .insn_retry(decode_retry),// set if branch_target_retry AND new inst_valid (always false in lab3)
  .insn_valid(decode_valid), 
    .insn(decode_insn), 

    .pc(decode_pc),

    .sign_ext(decode_sign_ext), 
    .src1(rs1_data),//decode_src1), 
    .src2(rs2_data),//decode_src2),
    .rd(decode_insn[11:7]),

    // From execute to register file (decode)
    // No need, RF always accepts writes input         dest_retry, 
    .dest_valid(dest_valid),
    .dest_retry(dest_retry),
    .dest_rd(dest_rd),
    .dest_long(dest_long),
    .dest_data(dest_data),
    .dest_clear(dest_clear),    

    // From execute to fetch
    .branch_target_retry(execute_retry), 
    .branch_target_valid(execute_valid),
    .branch_target(execute_pc),

    // From execute to dcache
    .dcache_req_addr(dcache_req_addr),
    .dcache_req_data(dcache_req_data),
    .dcache_req_op(dcache_req_op),
    .dcache_req_rd(dcache_req_rd),
    .dcache_req_valid(dcache_req_valid),
    .dcache_req_retry(dcache_req_retry)

  );

//from execute to decode
/*
fflop #(.Size(5+64))ff_pc_rd ( 
  .din({dest_rd_next, }), 
  .dinValid(decode_valid), 
  .dinRetry(decode_retry), 

  .q({dest_rd, }),
  .qValid(),
  .qRetry(dcache_req_retry),
  .*);
  */

  //flop_e #(.Bits(5))dregflop ( .clk(clk), .reset(reset), .we(decode_valid), .d(dest_rd_next), .q(dest_rd));

  endmodule

