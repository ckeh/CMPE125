
package myaluops;

  const logic DO_ADD = 4'b1010;
  const logic DO_SUB = 4'b1111;

endpackage

